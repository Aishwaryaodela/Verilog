module and_gate1(input a,b, output c);
endmodule
