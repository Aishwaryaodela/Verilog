module or_gate(input a,b , output c);
endmodule
